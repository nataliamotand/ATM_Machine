library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity atm is
    port (
        clk : in std_logic;
        reset : in std_logic;
    );
end atm;

architecture behavioral of atm is

begin

end behavioral;